module sync2

import time

pub fn thread_yield() {
	time.sleep_ms(0)
}