module sync2

fn C.GetCurrentThreadId() u32

fn C.SetThreadDescription() int

fn C._mm_pause()